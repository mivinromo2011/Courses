module downcounter_testbench();
reg clk, reset;
wire [3:0] counter;

down_counter dut(clk, reset, counter);
initial begin
    $monitor("%b,  %b,  %b",clk,reset,counter);
clk=0;
forever #5 clk=~clk;
end
initial begin
reset=1;
#20;
reset=0;
end
endmodule
